module shiftLeft(
    input  [31:0] A,
    input  [31:0] B,
    output [31:0] Result
);

reg [31:0] temp;
integer i;

always @(A or B)
begin
    temp = 32'b0;

    if (B < 32)
    begin
        for (i = B; i < 32; i = i + 1)
        begin
            temp[i] = A[i-B];
        end
    end
end

assign Result = temp;

endmodule
