`timescale 1ns/1ps
module tb_AND;

  reg  [31:0] A_and, B_and;
  wire [31:0] Result_and;

  AND dut (A_and, B_and, Result_and);

  initial begin
    A_and = 0;          B_and = 0;          #10;
    A_and = 32'hAAAA;   B_and = 32'h5555;   #10;
    A_and = 32'hFFFF;   B_and = 32'h0F0F;   #10;
    A_and = 32'hDEAD;   B_and = 32'hDEAD;   #10;
    $finish;
  end

endmodule